Lorem ipsum dolor sit amet, consectetur adipiscing elit. Cras eu felis magna. Lorem ipsum dolor sit amet, consectetur adipiscing elit. Etiam nec quam sed nisi tincidunt dictum ac eu nisi. Pellentesque habitant morbi tristique senectus et netus et malesuada fames ac turpis egestas. Ut malesuada, purus eu egestas lacinia, magna felis interdum urna, in rhoncus dolor nisl at augue. Interdum et malesuada fames ac ante ipsum primis in faucibus. In in nulla eget diam rutrum bibendum. Orci varius natoque penatibus et magnis dis parturient montes, nascetur ridiculus mus.

Sed tellus ipsum, vestibulum condimentum arcu at, pretium maximus nulla. Nam risus quam, sodales at elit id, fermentum vestibulum nisi. Etiam a sollicitudin diam, a feugiat ante. Morbi in luctus nisl, sed pulvinar leo. Cras auctor felis et pellentesque pellentesque. Nam vitae placerat sapien, quis sagittis dolor. Aenean lectus tortor, tempor in sollicitudin sollicitudin, vehicula iaculis ex. Cras tempor tellus quis consectetur porttitor. Integer at dui ex. Donec sem erat, cursus non lacus eu, auctor tempus neque. Proin ac tellus ac turpis hendrerit tempus.

Donec massa sem, feugiat vel arcu vel, ullamcorper malesuada ipsum. Suspendisse odio eros, auctor eu venenatis in, pharetra non odio. Class aptent taciti sociosqu ad litora torquent per conubia nostra, per inceptos himenaeos. Integer lobortis ut lectus sed eleifend. Nulla at odio non neque lacinia eleifend at eget libero. Suspendisse maximus sed dolor eget scelerisque. Nullam ut scelerisque justo. Class aptent taciti sociosqu ad litora torquent per conubia nostra, per inceptos himenaeos. Praesent vitae justo posuere, porttitor turpis vel, porttitor augue. Fusce vitae ante metus. Donec justo orci, condimentum vitae cursus at, consectetur quis ligula. Sed eu dolor vel diam vulputate tristique in non velit. Fusce pharetra ligula eget sapien pellentesque, nec pretium metus efficitur.

Nam et odio a velit tincidunt sollicitudin vitae non orci. Duis vehicula magna felis, vitae interdum quam tempor vitae. Aliquam eu lorem et massa commodo imperdiet. Curabitur mattis urna augue, a dictum massa scelerisque quis. Sed id arcu congue, hendrerit elit quis, egestas odio. Nullam eu lobortis sem. Sed dapibus tincidunt orci a luctus.

Nunc euismod, felis sit amet interdum iaculis, lorem ante vestibulum elit, id varius ligula augue quis ex. Vestibulum ante ipsum primis in faucibus orci luctus et ultrices posuere cubilia curae; Integer porttitor sem posuere pellentesque pharetra. Vestibulum ornare mauris sit amet sollicitudin molestie. Proin non faucibus dolor, vel venenatis ligula. Praesent tristique ipsum vel eros ornare, a sagittis elit imperdiet. Morbi elementum, enim sed interdum placerat, ipsum lacus vulputate dui, sodales pulvinar ex dolor in mi. Cras dapibus ex a tortor facilisis, sed vulputate nunc tincidunt. In posuere molestie porttitor. Vestibulum ante ipsum primis in faucibus orci luctus et ultrices posuere cubilia curae; Vestibulum aliquet arcu eget blandit tempus. Integer consectetur nunc nisi, at euismod nisi porta in. Curabitur in elit fringilla, ultrices nibh in, auctor nunc. Nam id nisi dapibus ex ornare sodales vitae a elit. Praesent sed velit at metus pharetra finibus nec quis libero.

Nullam in enim eget felis fringilla pulvinar et sed ipsum. Aliquam faucibus eros nec lectus maximus tincidunt. Nam vulputate ante vehicula mi commodo maximus. Mauris tellus libero, rhoncus in erat nec, sollicitudin lacinia ipsum. Pellentesque non congue erat. Etiam mattis est at bibendum tempor. Cras non nunc porta nunc elementum fermentum. Suspendisse sagittis ipsum et ex dictum porta. Cras a metus sed mauris lacinia condimentum sit amet eget erat. Nunc in sollicitudin lorem. Integer et justo finibus, pharetra arcu eget, tincidunt tortor. Quisque lectus nunc, lobortis et sagittis at, mollis sit amet nisi. Aliquam erat volutpat. Aenean lorem sem, varius eu mi in, egestas ultricies ipsum. Donec rutrum nibh et congue tempus. Quisque feugiat, libero nec sollicitudin laoreet, nulla ipsum placerat leo, quis ullamcorper tortor arcu eu odio.

Pellentesque et arcu nunc. In hac habitasse platea dictumst. In hac habitasse platea dictumst. Nam placerat hendrerit lacus vitae luctus. Etiam fringilla quam id molestie tempus. Nullam id ante dui. Fusce nec sagittis mi, eget fringilla dolor. Nullam sem nunc, eleifend eget luctus nec, efficitur et nulla. Nam faucibus massa sit amet lacinia aliquam.

Maecenas eu pharetra arcu. Nullam quis lorem sed ipsum hendrerit dictum et at metus. Aenean rhoncus tellus metus, quis varius velit viverra a. In tempus nisl ut maximus auctor. Phasellus sagittis diam turpis, non venenatis eros blandit ut. Phasellus elementum molestie risus, eget congue purus rutrum eget. Cras eu lorem eros. Praesent ac dui nibh. Etiam leo erat, tempor feugiat viverra quis, ullamcorper fringilla quam. Quisque vestibulum risus quis eros congue, nec ultrices erat consequat. Integer porta ex et ullamcorper maximus.

Nulla facilisi. Cras lobortis, nibh eget facilisis auctor, libero enim scelerisque odio, vel auctor libero mi in risus. Ut in finibus leo. Maecenas pellentesque laoreet turpis luctus lacinia. Maecenas vitae ex luctus, imperdiet augue egestas, posuere nisi. Morbi et mauris pulvinar, maximus augue at, tristique tortor. Donec lobortis hendrerit eleifend. Donec a enim vel quam rutrum congue ut quis nisl. Suspendisse hendrerit condimentum pellentesque. Aenean finibus risus nunc, ac suscipit massa tempor sed. Nunc lobortis commodo quam, id mollis quam pharetra quis. Donec sit amet nunc dolor.

Integer euismod suscipit ante id venenatis. Morbi vitae nulla molestie, euismod erat at, dapibus turpis. Sed condimentum felis nibh, et lacinia leo pretium vitae. Etiam sit amet elit a dui interdum sodales. Sed pharetra lacus quam, id ornare libero laoreet vitae. Aenean varius tellus at convallis dictum. Fusce interdum, mauris at convallis porta, est felis rhoncus enim, convallis commodo lorem libero non justo. Mauris congue volutpat sagittis.

Phasellus efficitur tincidunt nisl mattis venenatis. Nam at justo id turpis maximus interdum. Nulla ut convallis velit, sed sagittis sapien. Sed posuere lacinia orci eget fermentum. Donec pharetra massa eu tellus consequat, sed imperdiet justo suscipit. Aenean aliquet venenatis felis sed egestas. Fusce varius enim ut tincidunt varius. Donec at iaculis neque, eget tincidunt enim. Fusce posuere, lacus sit amet mollis ultricies, velit est congue purus, ut imperdiet massa purus vitae lectus. Aliquam facilisis nulla sit amet sem auctor, vel vulputate lorem scelerisque. In enim tellus, aliquam nec diam sit amet, convallis ullamcorper mi. Donec eget leo quis odio fringilla elementum.

Duis vitae fermentum nibh. Vestibulum non blandit nisl, eu congue ligula. Nulla ornare quam non mattis porttitor. Aliquam imperdiet dolor massa, sit amet semper velit aliquet at. Lorem ipsum dolor sit amet, consectetur adipiscing elit. Nam blandit sapien tellus, nec feugiat justo eleifend eu. Nulla ullamcorper sapien a aliquet tempus. Vestibulum vel pulvinar diam. Nam viverra ullamcorper erat id malesuada. Sed id ornare neque. Aliquam gravida consequat nibh euismod placerat. Donec placerat, tortor in finibus euismod, leo dolor laoreet lorem, tincidunt porta justo est at lorem. Sed auctor, augue non mattis finibus, urna sem mollis nisi, eu tristique turpis diam convallis elit. Aliquam non porttitor magna. Nam sollicitudin convallis tincidunt.

Curabitur dignissim interdum ex quis euismod. Duis posuere pharetra pharetra. Mauris malesuada mauris vel maximus convallis. Ut sodales lacinia malesuada. Suspendisse venenatis enim sit amet mattis maximus. Morbi finibus laoreet odio, sit amet facilisis tellus aliquam et. Proin posuere diam ligula, nec tincidunt purus rutrum at. Curabitur id congue massa. Ut malesuada condimentum enim id rhoncus.

Mauris erat lorem, porttitor eu nisi sed, rhoncus auctor erat. Morbi accumsan nisl non cursus scelerisque. Nulla facilisi. Pellentesque eu ante mollis mi semper tempus at sed velit. Donec sed maximus elit. Suspendisse non ex in nunc convallis rutrum. Aliquam non elit ipsum. Nullam vulputate ullamcorper velit. Ut ac magna lectus. Nullam placerat nulla in auctor elementum.

Sed eget lorem vitae justo iaculis consectetur. Donec id posuere justo. Ut maximus accumsan tellus eget aliquam. Nam eu accumsan purus. Etiam auctor risus nunc, in commodo enim eleifend volutpat. Praesent urna sapien, porttitor eget sem eu, sagittis iaculis lorem. Curabitur vitae semper augue. Aliquam sit amet ullamcorper tortor, vel sagittis odio.
